`include "subtracter/sub.v"
`include "subtracter/sub4.v"
module sub64( a, b, c, d, br);
input [63:0]a, b;
input c;
output [63:0]d;
output br;
wire [63:0]w;

sub4 s0(a[3:0],b[3:0],c,d[3:0],w[0]);
sub4 s1(a[7:4],b[7:4],w[0],d[7:4],w[1]);
sub4 s2(a[11:8],b[11:8],w[1],d[11:8],w[2]);
sub4 s3(a[15:12],b[15:12],w[2],d[15:12],w[3]);
sub4 s4(a[19:16],b[19:16],w[3],d[19:16],w[4]);
sub4 s5(a[23:20],b[23:20],w[4],d[23:20],w[5]);
sub4 s6(a[27:24],b[27:24],w[5],d[27:24],w[6]);
sub4 s7(a[31:28],b[31:28],w[6],d[31:28],w[7]);
sub4 s8(a[35:32],b[35:32],w[7],d[35:32],w[8]);
sub4 s9(a[39:36],b[39:36],w[8],d[39:36],w[9]);
sub4 s10(a[43:40],b[43:40],w[9],d[43:40],w[10]);
sub4 s11(a[47:44],b[47:44],w[10],d[47:44],w[11]);
sub4 s12(a[51:48],b[51:48],w[11],d[51:48],w[12]);
sub4 s13(a[55:52],b[55:52],w[12],d[55:52],w[13]);
sub4 s14(a[59:56],b[59:56],w[13],d[59:56],w[14]);
sub4 s15(a[63:60],b[63:60],w[14],d[63:60],br);

endmodule