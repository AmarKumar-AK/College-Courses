module example
(
 input x,
 input y,
 input z,
 output A,
 );

xor G1(A,x,y,z)

endmodule
